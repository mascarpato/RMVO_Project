library IEEE;
use IEEE.STD_LOGIC_1164.all;

package target is

type iu_config_type is record
	testboolean			:	boolean;
	testboolean2		:	boolean;
	testinteger			:	integer;
	data_memory_width	:	integer;
end record;

end target;

package body target is
end target;